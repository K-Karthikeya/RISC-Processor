// one-hot encoding for set_enable
module decoder_6_64(
  input [5:0] index,
  output [63:0] cacheline_meta	// cache line to be read from
);

// decoding the cache lines to be read from 
assign cacheline_meta = 	  (index == 0)	?	64'h1		:
                            (index == 1)	?	64'h2		:
                            (index == 2)	?	64'h4	    :
                            (index == 3)	?	64'h8	    :
                            (index == 4)	?	64'h10	    :
                            (index == 5)	?	64'h20	    :
                            (index == 6)	?	64'h40		:
                            (index == 7)	?	64'h80	    :
                            (index == 8)	?	64'h100	    :
                            (index == 9)	?	64'h200     :	
                            (index == 10)	?	64'h400     :
                            (index == 11)	?	64'h800     :
                            (index == 12)	?	64'h1000    :
                            (index == 13)	?	64'h2000    :
                            (index == 14)	?	64'h4000    :
                            (index == 15)   ?   64'h8000    :
                            (index == 16)   ?   64'h10000   :
                            (index == 17)   ?   64'h20000   :
                            (index == 18)   ?   64'h40000   :
                            (index == 19)   ?   64'h80000   :
                            (index == 20)   ?   64'h100000  :
                            (index == 21)   ?   64'h200000  :
                            (index == 22)   ?   64'h400000  :
                            (index == 23)   ?   64'h800000  :
                            (index == 24)   ?   64'h1000000 :
                            (index == 25)   ?   64'h2000000 :
                            (index == 26)   ?   64'h4000000 :
                            (index == 27)   ?   64'h8000000 :
                            (index == 28)   ?   64'h10000000    :
                            (index == 29)   ?   64'h20000000    :
                            (index == 30)   ?   64'h40000000    :
                            (index == 31)   ?   64'h80000000    :
                            (index == 32)   ?   64'h100000000   :
                            (index == 33)   ?   64'h200000000   :
                            (index == 34)   ?   64'h400000000   :   
                            (index == 35)   ?   64'h800000000   :
                            (index == 36)   ?   64'h1000000000  :
                            (index == 37)   ?   64'h2000000000  :
                            (index == 38)   ?   64'h4000000000  :
                            (index == 39)   ?   64'h8000000000  :
                            (index == 40)   ?   64'h10000000000 :
                            (index == 41)   ?   64'h20000000000 :
                            (index == 42)   ?   64'h40000000000 :
                            (index == 43)   ?   64'h80000000000 :
                            (index == 44)   ?   64'h100000000000    :
                            (index == 45)   ?   64'h200000000000    :
                            (index == 46)   ?   64'h400000000000    :
                            (index == 47)   ?   64'h800000000000    :
                            (index == 48)   ?   64'h1000000000000   :
                            (index == 49)   ?   64'h2000000000000   :
                            (index == 50)   ?   64'h4000000000000   :
                            (index == 51)   ?   64'h8000000000000   :
                            (index == 52)   ?   64'h10000000000000  :
                            (index == 53)   ?   64'h20000000000000  :
                            (index == 54)   ?   64'h40000000000000  :
                            (index == 55)   ?   64'h80000000000000  :
                            (index == 56)   ?   64'h100000000000000 :
                            (index == 57)   ?   64'h200000000000000 :
                            (index == 58)   ?   64'h400000000000000 :
                            (index == 59)   ?   64'h800000000000000 :
                            (index == 60)   ?   64'h1000000000000000    :
                            (index == 61)   ?   64'h2000000000000000    :
                            (index == 62)   ?   64'h4000000000000000    :
                                                64'h8000000000000000;


endmodule		// decoder